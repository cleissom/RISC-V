use std.textio.all;

package constants is
	constant data_width : integer := 32;
	constant dmemory_size : integer := 32;
	constant imemory_width : integer := 10;
	constant dmemory_width : integer := 10;
	constant memory_file : string := "code.txt";
end package constants;

package body constants is
end package body constants;
