use std.textio.all;

package constants is
	constant data_width : integer := 32;
	constant dmemory_size : integer := 32;
end package constants;

package body constants is
end package body constants;
